// soc_ethond.v

// Generated using ACDS version 14.0 200 at 2015.11.25.12:59:52

`timescale 1 ps / 1 ps
module soc_ethond (
		output wire [14:0] memory_mem_a,                     //        memory.mem_a
		output wire [2:0]  memory_mem_ba,                    //              .mem_ba
		output wire        memory_mem_ck,                    //              .mem_ck
		output wire        memory_mem_ck_n,                  //              .mem_ck_n
		output wire        memory_mem_cke,                   //              .mem_cke
		output wire        memory_mem_cs_n,                  //              .mem_cs_n
		output wire        memory_mem_ras_n,                 //              .mem_ras_n
		output wire        memory_mem_cas_n,                 //              .mem_cas_n
		output wire        memory_mem_we_n,                  //              .mem_we_n
		output wire        memory_mem_reset_n,               //              .mem_reset_n
		inout  wire [31:0] memory_mem_dq,                    //              .mem_dq
		inout  wire [3:0]  memory_mem_dqs,                   //              .mem_dqs
		inout  wire [3:0]  memory_mem_dqs_n,                 //              .mem_dqs_n
		output wire        memory_mem_odt,                   //              .mem_odt
		output wire [3:0]  memory_mem_dm,                    //              .mem_dm
		input  wire        memory_oct_rzqin,                 //              .oct_rzqin
		output wire        hps_io_hps_io_emac1_inst_TX_CLK,  //        hps_io.hps_io_emac1_inst_TX_CLK
		output wire        hps_io_hps_io_emac1_inst_TXD0,    //              .hps_io_emac1_inst_TXD0
		output wire        hps_io_hps_io_emac1_inst_TXD1,    //              .hps_io_emac1_inst_TXD1
		output wire        hps_io_hps_io_emac1_inst_TXD2,    //              .hps_io_emac1_inst_TXD2
		output wire        hps_io_hps_io_emac1_inst_TXD3,    //              .hps_io_emac1_inst_TXD3
		input  wire        hps_io_hps_io_emac1_inst_RXD0,    //              .hps_io_emac1_inst_RXD0
		inout  wire        hps_io_hps_io_emac1_inst_MDIO,    //              .hps_io_emac1_inst_MDIO
		output wire        hps_io_hps_io_emac1_inst_MDC,     //              .hps_io_emac1_inst_MDC
		input  wire        hps_io_hps_io_emac1_inst_RX_CTL,  //              .hps_io_emac1_inst_RX_CTL
		output wire        hps_io_hps_io_emac1_inst_TX_CTL,  //              .hps_io_emac1_inst_TX_CTL
		input  wire        hps_io_hps_io_emac1_inst_RX_CLK,  //              .hps_io_emac1_inst_RX_CLK
		input  wire        hps_io_hps_io_emac1_inst_RXD1,    //              .hps_io_emac1_inst_RXD1
		input  wire        hps_io_hps_io_emac1_inst_RXD2,    //              .hps_io_emac1_inst_RXD2
		input  wire        hps_io_hps_io_emac1_inst_RXD3,    //              .hps_io_emac1_inst_RXD3
		inout  wire        hps_io_hps_io_qspi_inst_IO0,      //              .hps_io_qspi_inst_IO0
		inout  wire        hps_io_hps_io_qspi_inst_IO1,      //              .hps_io_qspi_inst_IO1
		inout  wire        hps_io_hps_io_qspi_inst_IO2,      //              .hps_io_qspi_inst_IO2
		inout  wire        hps_io_hps_io_qspi_inst_IO3,      //              .hps_io_qspi_inst_IO3
		output wire        hps_io_hps_io_qspi_inst_SS0,      //              .hps_io_qspi_inst_SS0
		output wire        hps_io_hps_io_qspi_inst_CLK,      //              .hps_io_qspi_inst_CLK
		inout  wire        hps_io_hps_io_sdio_inst_CMD,      //              .hps_io_sdio_inst_CMD
		inout  wire        hps_io_hps_io_sdio_inst_D0,       //              .hps_io_sdio_inst_D0
		inout  wire        hps_io_hps_io_sdio_inst_D1,       //              .hps_io_sdio_inst_D1
		output wire        hps_io_hps_io_sdio_inst_CLK,      //              .hps_io_sdio_inst_CLK
		inout  wire        hps_io_hps_io_sdio_inst_D2,       //              .hps_io_sdio_inst_D2
		inout  wire        hps_io_hps_io_sdio_inst_D3,       //              .hps_io_sdio_inst_D3
		inout  wire        hps_io_hps_io_usb1_inst_D0,       //              .hps_io_usb1_inst_D0
		inout  wire        hps_io_hps_io_usb1_inst_D1,       //              .hps_io_usb1_inst_D1
		inout  wire        hps_io_hps_io_usb1_inst_D2,       //              .hps_io_usb1_inst_D2
		inout  wire        hps_io_hps_io_usb1_inst_D3,       //              .hps_io_usb1_inst_D3
		inout  wire        hps_io_hps_io_usb1_inst_D4,       //              .hps_io_usb1_inst_D4
		inout  wire        hps_io_hps_io_usb1_inst_D5,       //              .hps_io_usb1_inst_D5
		inout  wire        hps_io_hps_io_usb1_inst_D6,       //              .hps_io_usb1_inst_D6
		inout  wire        hps_io_hps_io_usb1_inst_D7,       //              .hps_io_usb1_inst_D7
		input  wire        hps_io_hps_io_usb1_inst_CLK,      //              .hps_io_usb1_inst_CLK
		output wire        hps_io_hps_io_usb1_inst_STP,      //              .hps_io_usb1_inst_STP
		input  wire        hps_io_hps_io_usb1_inst_DIR,      //              .hps_io_usb1_inst_DIR
		input  wire        hps_io_hps_io_usb1_inst_NXT,      //              .hps_io_usb1_inst_NXT
		input  wire        hps_io_hps_io_uart0_inst_RX,      //              .hps_io_uart0_inst_RX
		output wire        hps_io_hps_io_uart0_inst_TX,      //              .hps_io_uart0_inst_TX
		inout  wire        hps_io_hps_io_i2c0_inst_SDA,      //              .hps_io_i2c0_inst_SDA
		inout  wire        hps_io_hps_io_i2c0_inst_SCL,      //              .hps_io_i2c0_inst_SCL
		inout  wire        hps_io_hps_io_gpio_inst_GPIO09,   //              .hps_io_gpio_inst_GPIO09
		inout  wire        hps_io_hps_io_gpio_inst_GPIO37,   //              .hps_io_gpio_inst_GPIO37
		inout  wire        hps_io_hps_io_gpio_inst_GPIO44,   //              .hps_io_gpio_inst_GPIO44
		inout  wire        hps_io_hps_io_gpio_inst_GPIO48,   //              .hps_io_gpio_inst_GPIO48
		inout  wire        hps_io_hps_io_gpio_inst_GPIO52,   //              .hps_io_gpio_inst_GPIO52
		inout  wire        hps_io_hps_io_gpio_inst_GPIO65,   //              .hps_io_gpio_inst_GPIO65
		inout  wire        hps_io_hps_io_gpio_inst_LOANIO58, //              .hps_io_gpio_inst_LOANIO58
		input  wire        sys_clk_clk,                      //       sys_clk.clk
		output wire        sys_rst_reset,                    //       sys_rst.reset
		output wire [66:0] hps_loan_io_in,                   //   hps_loan_io.in
		input  wire [66:0] hps_loan_io_out,                  //              .out
		input  wire [66:0] hps_loan_io_oe,                   //              .oe
		input  wire [31:0] irq0_irq,                         //          irq0.irq
		input  wire [31:0] irq1_irq,                         //          irq1.irq
		input  wire        netdma_csr0_waitrequest,          //   netdma_csr0.waitrequest
		input  wire [31:0] netdma_csr0_readdata,             //              .readdata
		input  wire        netdma_csr0_readdatavalid,        //              .readdatavalid
		output wire [0:0]  netdma_csr0_burstcount,           //              .burstcount
		output wire [31:0] netdma_csr0_writedata,            //              .writedata
		output wire [12:0] netdma_csr0_address,              //              .address
		output wire        netdma_csr0_write,                //              .write
		output wire        netdma_csr0_read,                 //              .read
		output wire [3:0]  netdma_csr0_byteenable,           //              .byteenable
		output wire        netdma_csr0_debugaccess,          //              .debugaccess
		input  wire        netdma_csr1_waitrequest,          //   netdma_csr1.waitrequest
		input  wire [31:0] netdma_csr1_readdata,             //              .readdata
		input  wire        netdma_csr1_readdatavalid,        //              .readdatavalid
		output wire [0:0]  netdma_csr1_burstcount,           //              .burstcount
		output wire [31:0] netdma_csr1_writedata,            //              .writedata
		output wire [12:0] netdma_csr1_address,              //              .address
		output wire        netdma_csr1_write,                //              .write
		output wire        netdma_csr1_read,                 //              .read
		output wire [3:0]  netdma_csr1_byteenable,           //              .byteenable
		output wire        netdma_csr1_debugaccess,          //              .debugaccess
		output wire        netdma_write0_waitrequest,        // netdma_write0.waitrequest
		output wire [63:0] netdma_write0_readdata,           //              .readdata
		output wire        netdma_write0_readdatavalid,      //              .readdatavalid
		input  wire [0:0]  netdma_write0_burstcount,         //              .burstcount
		input  wire [63:0] netdma_write0_writedata,          //              .writedata
		input  wire [31:0] netdma_write0_address,            //              .address
		input  wire        netdma_write0_write,              //              .write
		input  wire        netdma_write0_read,               //              .read
		input  wire [7:0]  netdma_write0_byteenable,         //              .byteenable
		input  wire        netdma_write0_debugaccess,        //              .debugaccess
		output wire        netdma_write1_waitrequest,        // netdma_write1.waitrequest
		output wire [63:0] netdma_write1_readdata,           //              .readdata
		output wire        netdma_write1_readdatavalid,      //              .readdatavalid
		input  wire [0:0]  netdma_write1_burstcount,         //              .burstcount
		input  wire [63:0] netdma_write1_writedata,          //              .writedata
		input  wire [31:0] netdma_write1_address,            //              .address
		input  wire        netdma_write1_write,              //              .write
		input  wire        netdma_write1_read,               //              .read
		input  wire [7:0]  netdma_write1_byteenable,         //              .byteenable
		input  wire        netdma_write1_debugaccess,        //              .debugaccess
		output wire        netdma_read0_waitrequest,         //  netdma_read0.waitrequest
		output wire [63:0] netdma_read0_readdata,            //              .readdata
		output wire        netdma_read0_readdatavalid,       //              .readdatavalid
		input  wire [0:0]  netdma_read0_burstcount,          //              .burstcount
		input  wire [63:0] netdma_read0_writedata,           //              .writedata
		input  wire [31:0] netdma_read0_address,             //              .address
		input  wire        netdma_read0_write,               //              .write
		input  wire        netdma_read0_read,                //              .read
		input  wire [7:0]  netdma_read0_byteenable,          //              .byteenable
		input  wire        netdma_read0_debugaccess,         //              .debugaccess
		output wire        netdma_read1_waitrequest,         //  netdma_read1.waitrequest
		output wire [63:0] netdma_read1_readdata,            //              .readdata
		output wire        netdma_read1_readdatavalid,       //              .readdatavalid
		input  wire [0:0]  netdma_read1_burstcount,          //              .burstcount
		input  wire [63:0] netdma_read1_writedata,           //              .writedata
		input  wire [31:0] netdma_read1_address,             //              .address
		input  wire        netdma_read1_write,               //              .write
		input  wire        netdma_read1_read,                //              .read
		input  wire [7:0]  netdma_read1_byteenable,          //              .byteenable
		input  wire        netdma_read1_debugaccess,         //              .debugaccess
		input  wire        csr_waitrequest,                  //           csr.waitrequest
		input  wire [31:0] csr_readdata,                     //              .readdata
		input  wire        csr_readdatavalid,                //              .readdatavalid
		output wire [0:0]  csr_burstcount,                   //              .burstcount
		output wire [31:0] csr_writedata,                    //              .writedata
		output wire [12:0] csr_address,                      //              .address
		output wire        csr_write,                        //              .write
		output wire        csr_read,                         //              .read
		output wire [3:0]  csr_byteenable,                   //              .byteenable
		output wire        csr_debugaccess                   //              .debugaccess
	);

	wire         hps_0_h2f_axi_master_awvalid;                   // hps_0:h2f_AWVALID -> mm_interconnect_0:hps_0_h2f_axi_master_awvalid
	wire   [2:0] hps_0_h2f_axi_master_arsize;                    // hps_0:h2f_ARSIZE -> mm_interconnect_0:hps_0_h2f_axi_master_arsize
	wire   [1:0] hps_0_h2f_axi_master_arlock;                    // hps_0:h2f_ARLOCK -> mm_interconnect_0:hps_0_h2f_axi_master_arlock
	wire   [3:0] hps_0_h2f_axi_master_awcache;                   // hps_0:h2f_AWCACHE -> mm_interconnect_0:hps_0_h2f_axi_master_awcache
	wire         hps_0_h2f_axi_master_arready;                   // mm_interconnect_0:hps_0_h2f_axi_master_arready -> hps_0:h2f_ARREADY
	wire  [11:0] hps_0_h2f_axi_master_arid;                      // hps_0:h2f_ARID -> mm_interconnect_0:hps_0_h2f_axi_master_arid
	wire         hps_0_h2f_axi_master_rready;                    // hps_0:h2f_RREADY -> mm_interconnect_0:hps_0_h2f_axi_master_rready
	wire         hps_0_h2f_axi_master_bready;                    // hps_0:h2f_BREADY -> mm_interconnect_0:hps_0_h2f_axi_master_bready
	wire   [2:0] hps_0_h2f_axi_master_awsize;                    // hps_0:h2f_AWSIZE -> mm_interconnect_0:hps_0_h2f_axi_master_awsize
	wire   [2:0] hps_0_h2f_axi_master_awprot;                    // hps_0:h2f_AWPROT -> mm_interconnect_0:hps_0_h2f_axi_master_awprot
	wire         hps_0_h2f_axi_master_arvalid;                   // hps_0:h2f_ARVALID -> mm_interconnect_0:hps_0_h2f_axi_master_arvalid
	wire   [2:0] hps_0_h2f_axi_master_arprot;                    // hps_0:h2f_ARPROT -> mm_interconnect_0:hps_0_h2f_axi_master_arprot
	wire  [11:0] hps_0_h2f_axi_master_bid;                       // mm_interconnect_0:hps_0_h2f_axi_master_bid -> hps_0:h2f_BID
	wire   [3:0] hps_0_h2f_axi_master_arlen;                     // hps_0:h2f_ARLEN -> mm_interconnect_0:hps_0_h2f_axi_master_arlen
	wire         hps_0_h2f_axi_master_awready;                   // mm_interconnect_0:hps_0_h2f_axi_master_awready -> hps_0:h2f_AWREADY
	wire  [11:0] hps_0_h2f_axi_master_awid;                      // hps_0:h2f_AWID -> mm_interconnect_0:hps_0_h2f_axi_master_awid
	wire         hps_0_h2f_axi_master_bvalid;                    // mm_interconnect_0:hps_0_h2f_axi_master_bvalid -> hps_0:h2f_BVALID
	wire  [11:0] hps_0_h2f_axi_master_wid;                       // hps_0:h2f_WID -> mm_interconnect_0:hps_0_h2f_axi_master_wid
	wire   [1:0] hps_0_h2f_axi_master_awlock;                    // hps_0:h2f_AWLOCK -> mm_interconnect_0:hps_0_h2f_axi_master_awlock
	wire   [1:0] hps_0_h2f_axi_master_awburst;                   // hps_0:h2f_AWBURST -> mm_interconnect_0:hps_0_h2f_axi_master_awburst
	wire   [1:0] hps_0_h2f_axi_master_bresp;                     // mm_interconnect_0:hps_0_h2f_axi_master_bresp -> hps_0:h2f_BRESP
	wire   [3:0] hps_0_h2f_axi_master_wstrb;                     // hps_0:h2f_WSTRB -> mm_interconnect_0:hps_0_h2f_axi_master_wstrb
	wire         hps_0_h2f_axi_master_rvalid;                    // mm_interconnect_0:hps_0_h2f_axi_master_rvalid -> hps_0:h2f_RVALID
	wire  [31:0] hps_0_h2f_axi_master_wdata;                     // hps_0:h2f_WDATA -> mm_interconnect_0:hps_0_h2f_axi_master_wdata
	wire         hps_0_h2f_axi_master_wready;                    // mm_interconnect_0:hps_0_h2f_axi_master_wready -> hps_0:h2f_WREADY
	wire   [1:0] hps_0_h2f_axi_master_arburst;                   // hps_0:h2f_ARBURST -> mm_interconnect_0:hps_0_h2f_axi_master_arburst
	wire  [31:0] hps_0_h2f_axi_master_rdata;                     // mm_interconnect_0:hps_0_h2f_axi_master_rdata -> hps_0:h2f_RDATA
	wire  [29:0] hps_0_h2f_axi_master_araddr;                    // hps_0:h2f_ARADDR -> mm_interconnect_0:hps_0_h2f_axi_master_araddr
	wire   [3:0] hps_0_h2f_axi_master_arcache;                   // hps_0:h2f_ARCACHE -> mm_interconnect_0:hps_0_h2f_axi_master_arcache
	wire   [3:0] hps_0_h2f_axi_master_awlen;                     // hps_0:h2f_AWLEN -> mm_interconnect_0:hps_0_h2f_axi_master_awlen
	wire  [29:0] hps_0_h2f_axi_master_awaddr;                    // hps_0:h2f_AWADDR -> mm_interconnect_0:hps_0_h2f_axi_master_awaddr
	wire  [11:0] hps_0_h2f_axi_master_rid;                       // mm_interconnect_0:hps_0_h2f_axi_master_rid -> hps_0:h2f_RID
	wire         hps_0_h2f_axi_master_wvalid;                    // hps_0:h2f_WVALID -> mm_interconnect_0:hps_0_h2f_axi_master_wvalid
	wire   [1:0] hps_0_h2f_axi_master_rresp;                     // mm_interconnect_0:hps_0_h2f_axi_master_rresp -> hps_0:h2f_RRESP
	wire         hps_0_h2f_axi_master_wlast;                     // hps_0:h2f_WLAST -> mm_interconnect_0:hps_0_h2f_axi_master_wlast
	wire         hps_0_h2f_axi_master_rlast;                     // mm_interconnect_0:hps_0_h2f_axi_master_rlast -> hps_0:h2f_RLAST
	wire         mm_interconnect_0_mm_bridge_5_s0_waitrequest;   // mm_bridge_5:s0_waitrequest -> mm_interconnect_0:mm_bridge_5_s0_waitrequest
	wire   [0:0] mm_interconnect_0_mm_bridge_5_s0_burstcount;    // mm_interconnect_0:mm_bridge_5_s0_burstcount -> mm_bridge_5:s0_burstcount
	wire  [31:0] mm_interconnect_0_mm_bridge_5_s0_writedata;     // mm_interconnect_0:mm_bridge_5_s0_writedata -> mm_bridge_5:s0_writedata
	wire  [12:0] mm_interconnect_0_mm_bridge_5_s0_address;       // mm_interconnect_0:mm_bridge_5_s0_address -> mm_bridge_5:s0_address
	wire         mm_interconnect_0_mm_bridge_5_s0_write;         // mm_interconnect_0:mm_bridge_5_s0_write -> mm_bridge_5:s0_write
	wire         mm_interconnect_0_mm_bridge_5_s0_read;          // mm_interconnect_0:mm_bridge_5_s0_read -> mm_bridge_5:s0_read
	wire  [31:0] mm_interconnect_0_mm_bridge_5_s0_readdata;      // mm_bridge_5:s0_readdata -> mm_interconnect_0:mm_bridge_5_s0_readdata
	wire         mm_interconnect_0_mm_bridge_5_s0_debugaccess;   // mm_interconnect_0:mm_bridge_5_s0_debugaccess -> mm_bridge_5:s0_debugaccess
	wire         mm_interconnect_0_mm_bridge_5_s0_readdatavalid; // mm_bridge_5:s0_readdatavalid -> mm_interconnect_0:mm_bridge_5_s0_readdatavalid
	wire   [3:0] mm_interconnect_0_mm_bridge_5_s0_byteenable;    // mm_interconnect_0:mm_bridge_5_s0_byteenable -> mm_bridge_5:s0_byteenable
	wire         mm_interconnect_0_mm_bridge_6_s0_waitrequest;   // mm_bridge_6:s0_waitrequest -> mm_interconnect_0:mm_bridge_6_s0_waitrequest
	wire   [0:0] mm_interconnect_0_mm_bridge_6_s0_burstcount;    // mm_interconnect_0:mm_bridge_6_s0_burstcount -> mm_bridge_6:s0_burstcount
	wire  [31:0] mm_interconnect_0_mm_bridge_6_s0_writedata;     // mm_interconnect_0:mm_bridge_6_s0_writedata -> mm_bridge_6:s0_writedata
	wire  [12:0] mm_interconnect_0_mm_bridge_6_s0_address;       // mm_interconnect_0:mm_bridge_6_s0_address -> mm_bridge_6:s0_address
	wire         mm_interconnect_0_mm_bridge_6_s0_write;         // mm_interconnect_0:mm_bridge_6_s0_write -> mm_bridge_6:s0_write
	wire         mm_interconnect_0_mm_bridge_6_s0_read;          // mm_interconnect_0:mm_bridge_6_s0_read -> mm_bridge_6:s0_read
	wire  [31:0] mm_interconnect_0_mm_bridge_6_s0_readdata;      // mm_bridge_6:s0_readdata -> mm_interconnect_0:mm_bridge_6_s0_readdata
	wire         mm_interconnect_0_mm_bridge_6_s0_debugaccess;   // mm_interconnect_0:mm_bridge_6_s0_debugaccess -> mm_bridge_6:s0_debugaccess
	wire         mm_interconnect_0_mm_bridge_6_s0_readdatavalid; // mm_bridge_6:s0_readdatavalid -> mm_interconnect_0:mm_bridge_6_s0_readdatavalid
	wire   [3:0] mm_interconnect_0_mm_bridge_6_s0_byteenable;    // mm_interconnect_0:mm_bridge_6_s0_byteenable -> mm_bridge_6:s0_byteenable
	wire         mm_interconnect_0_mm_bridge_0_s0_waitrequest;   // mm_bridge_0:s0_waitrequest -> mm_interconnect_0:mm_bridge_0_s0_waitrequest
	wire   [0:0] mm_interconnect_0_mm_bridge_0_s0_burstcount;    // mm_interconnect_0:mm_bridge_0_s0_burstcount -> mm_bridge_0:s0_burstcount
	wire  [31:0] mm_interconnect_0_mm_bridge_0_s0_writedata;     // mm_interconnect_0:mm_bridge_0_s0_writedata -> mm_bridge_0:s0_writedata
	wire  [12:0] mm_interconnect_0_mm_bridge_0_s0_address;       // mm_interconnect_0:mm_bridge_0_s0_address -> mm_bridge_0:s0_address
	wire         mm_interconnect_0_mm_bridge_0_s0_write;         // mm_interconnect_0:mm_bridge_0_s0_write -> mm_bridge_0:s0_write
	wire         mm_interconnect_0_mm_bridge_0_s0_read;          // mm_interconnect_0:mm_bridge_0_s0_read -> mm_bridge_0:s0_read
	wire  [31:0] mm_interconnect_0_mm_bridge_0_s0_readdata;      // mm_bridge_0:s0_readdata -> mm_interconnect_0:mm_bridge_0_s0_readdata
	wire         mm_interconnect_0_mm_bridge_0_s0_debugaccess;   // mm_interconnect_0:mm_bridge_0_s0_debugaccess -> mm_bridge_0:s0_debugaccess
	wire         mm_interconnect_0_mm_bridge_0_s0_readdatavalid; // mm_bridge_0:s0_readdatavalid -> mm_interconnect_0:mm_bridge_0_s0_readdatavalid
	wire   [3:0] mm_interconnect_0_mm_bridge_0_s0_byteenable;    // mm_interconnect_0:mm_bridge_0_s0_byteenable -> mm_bridge_0:s0_byteenable
	wire   [0:0] mm_bridge_1_m0_burstcount;                      // mm_bridge_1:m0_burstcount -> mm_interconnect_1:mm_bridge_1_m0_burstcount
	wire         mm_bridge_1_m0_waitrequest;                     // mm_interconnect_1:mm_bridge_1_m0_waitrequest -> mm_bridge_1:m0_waitrequest
	wire  [31:0] mm_bridge_1_m0_address;                         // mm_bridge_1:m0_address -> mm_interconnect_1:mm_bridge_1_m0_address
	wire  [63:0] mm_bridge_1_m0_writedata;                       // mm_bridge_1:m0_writedata -> mm_interconnect_1:mm_bridge_1_m0_writedata
	wire         mm_bridge_1_m0_write;                           // mm_bridge_1:m0_write -> mm_interconnect_1:mm_bridge_1_m0_write
	wire         mm_bridge_1_m0_read;                            // mm_bridge_1:m0_read -> mm_interconnect_1:mm_bridge_1_m0_read
	wire  [63:0] mm_bridge_1_m0_readdata;                        // mm_interconnect_1:mm_bridge_1_m0_readdata -> mm_bridge_1:m0_readdata
	wire         mm_bridge_1_m0_debugaccess;                     // mm_bridge_1:m0_debugaccess -> mm_interconnect_1:mm_bridge_1_m0_debugaccess
	wire   [7:0] mm_bridge_1_m0_byteenable;                      // mm_bridge_1:m0_byteenable -> mm_interconnect_1:mm_bridge_1_m0_byteenable
	wire         mm_bridge_1_m0_readdatavalid;                   // mm_interconnect_1:mm_bridge_1_m0_readdatavalid -> mm_bridge_1:m0_readdatavalid
	wire   [0:0] mm_bridge_3_m0_burstcount;                      // mm_bridge_3:m0_burstcount -> mm_interconnect_1:mm_bridge_3_m0_burstcount
	wire         mm_bridge_3_m0_waitrequest;                     // mm_interconnect_1:mm_bridge_3_m0_waitrequest -> mm_bridge_3:m0_waitrequest
	wire  [31:0] mm_bridge_3_m0_address;                         // mm_bridge_3:m0_address -> mm_interconnect_1:mm_bridge_3_m0_address
	wire  [63:0] mm_bridge_3_m0_writedata;                       // mm_bridge_3:m0_writedata -> mm_interconnect_1:mm_bridge_3_m0_writedata
	wire         mm_bridge_3_m0_write;                           // mm_bridge_3:m0_write -> mm_interconnect_1:mm_bridge_3_m0_write
	wire         mm_bridge_3_m0_read;                            // mm_bridge_3:m0_read -> mm_interconnect_1:mm_bridge_3_m0_read
	wire  [63:0] mm_bridge_3_m0_readdata;                        // mm_interconnect_1:mm_bridge_3_m0_readdata -> mm_bridge_3:m0_readdata
	wire         mm_bridge_3_m0_debugaccess;                     // mm_bridge_3:m0_debugaccess -> mm_interconnect_1:mm_bridge_3_m0_debugaccess
	wire   [7:0] mm_bridge_3_m0_byteenable;                      // mm_bridge_3:m0_byteenable -> mm_interconnect_1:mm_bridge_3_m0_byteenable
	wire         mm_bridge_3_m0_readdatavalid;                   // mm_interconnect_1:mm_bridge_3_m0_readdatavalid -> mm_bridge_3:m0_readdatavalid
	wire   [0:0] mm_bridge_4_m0_burstcount;                      // mm_bridge_4:m0_burstcount -> mm_interconnect_1:mm_bridge_4_m0_burstcount
	wire         mm_bridge_4_m0_waitrequest;                     // mm_interconnect_1:mm_bridge_4_m0_waitrequest -> mm_bridge_4:m0_waitrequest
	wire  [31:0] mm_bridge_4_m0_address;                         // mm_bridge_4:m0_address -> mm_interconnect_1:mm_bridge_4_m0_address
	wire  [63:0] mm_bridge_4_m0_writedata;                       // mm_bridge_4:m0_writedata -> mm_interconnect_1:mm_bridge_4_m0_writedata
	wire         mm_bridge_4_m0_write;                           // mm_bridge_4:m0_write -> mm_interconnect_1:mm_bridge_4_m0_write
	wire         mm_bridge_4_m0_read;                            // mm_bridge_4:m0_read -> mm_interconnect_1:mm_bridge_4_m0_read
	wire  [63:0] mm_bridge_4_m0_readdata;                        // mm_interconnect_1:mm_bridge_4_m0_readdata -> mm_bridge_4:m0_readdata
	wire         mm_bridge_4_m0_debugaccess;                     // mm_bridge_4:m0_debugaccess -> mm_interconnect_1:mm_bridge_4_m0_debugaccess
	wire   [7:0] mm_bridge_4_m0_byteenable;                      // mm_bridge_4:m0_byteenable -> mm_interconnect_1:mm_bridge_4_m0_byteenable
	wire         mm_bridge_4_m0_readdatavalid;                   // mm_interconnect_1:mm_bridge_4_m0_readdatavalid -> mm_bridge_4:m0_readdatavalid
	wire   [0:0] mm_bridge_2_m0_burstcount;                      // mm_bridge_2:m0_burstcount -> mm_interconnect_1:mm_bridge_2_m0_burstcount
	wire         mm_bridge_2_m0_waitrequest;                     // mm_interconnect_1:mm_bridge_2_m0_waitrequest -> mm_bridge_2:m0_waitrequest
	wire  [31:0] mm_bridge_2_m0_address;                         // mm_bridge_2:m0_address -> mm_interconnect_1:mm_bridge_2_m0_address
	wire  [63:0] mm_bridge_2_m0_writedata;                       // mm_bridge_2:m0_writedata -> mm_interconnect_1:mm_bridge_2_m0_writedata
	wire         mm_bridge_2_m0_write;                           // mm_bridge_2:m0_write -> mm_interconnect_1:mm_bridge_2_m0_write
	wire         mm_bridge_2_m0_read;                            // mm_bridge_2:m0_read -> mm_interconnect_1:mm_bridge_2_m0_read
	wire  [63:0] mm_bridge_2_m0_readdata;                        // mm_interconnect_1:mm_bridge_2_m0_readdata -> mm_bridge_2:m0_readdata
	wire         mm_bridge_2_m0_debugaccess;                     // mm_bridge_2:m0_debugaccess -> mm_interconnect_1:mm_bridge_2_m0_debugaccess
	wire   [7:0] mm_bridge_2_m0_byteenable;                      // mm_bridge_2:m0_byteenable -> mm_interconnect_1:mm_bridge_2_m0_byteenable
	wire         mm_bridge_2_m0_readdatavalid;                   // mm_interconnect_1:mm_bridge_2_m0_readdatavalid -> mm_bridge_2:m0_readdatavalid
	wire         mm_interconnect_1_hps_0_f2h_axi_slave_awvalid;  // mm_interconnect_1:hps_0_f2h_axi_slave_awvalid -> hps_0:f2h_AWVALID
	wire   [2:0] mm_interconnect_1_hps_0_f2h_axi_slave_arsize;   // mm_interconnect_1:hps_0_f2h_axi_slave_arsize -> hps_0:f2h_ARSIZE
	wire   [1:0] mm_interconnect_1_hps_0_f2h_axi_slave_arlock;   // mm_interconnect_1:hps_0_f2h_axi_slave_arlock -> hps_0:f2h_ARLOCK
	wire   [3:0] mm_interconnect_1_hps_0_f2h_axi_slave_awcache;  // mm_interconnect_1:hps_0_f2h_axi_slave_awcache -> hps_0:f2h_AWCACHE
	wire         mm_interconnect_1_hps_0_f2h_axi_slave_arready;  // hps_0:f2h_ARREADY -> mm_interconnect_1:hps_0_f2h_axi_slave_arready
	wire   [7:0] mm_interconnect_1_hps_0_f2h_axi_slave_arid;     // mm_interconnect_1:hps_0_f2h_axi_slave_arid -> hps_0:f2h_ARID
	wire         mm_interconnect_1_hps_0_f2h_axi_slave_rready;   // mm_interconnect_1:hps_0_f2h_axi_slave_rready -> hps_0:f2h_RREADY
	wire         mm_interconnect_1_hps_0_f2h_axi_slave_bready;   // mm_interconnect_1:hps_0_f2h_axi_slave_bready -> hps_0:f2h_BREADY
	wire   [2:0] mm_interconnect_1_hps_0_f2h_axi_slave_awsize;   // mm_interconnect_1:hps_0_f2h_axi_slave_awsize -> hps_0:f2h_AWSIZE
	wire   [2:0] mm_interconnect_1_hps_0_f2h_axi_slave_awprot;   // mm_interconnect_1:hps_0_f2h_axi_slave_awprot -> hps_0:f2h_AWPROT
	wire         mm_interconnect_1_hps_0_f2h_axi_slave_arvalid;  // mm_interconnect_1:hps_0_f2h_axi_slave_arvalid -> hps_0:f2h_ARVALID
	wire   [2:0] mm_interconnect_1_hps_0_f2h_axi_slave_arprot;   // mm_interconnect_1:hps_0_f2h_axi_slave_arprot -> hps_0:f2h_ARPROT
	wire   [7:0] mm_interconnect_1_hps_0_f2h_axi_slave_bid;      // hps_0:f2h_BID -> mm_interconnect_1:hps_0_f2h_axi_slave_bid
	wire   [3:0] mm_interconnect_1_hps_0_f2h_axi_slave_arlen;    // mm_interconnect_1:hps_0_f2h_axi_slave_arlen -> hps_0:f2h_ARLEN
	wire         mm_interconnect_1_hps_0_f2h_axi_slave_awready;  // hps_0:f2h_AWREADY -> mm_interconnect_1:hps_0_f2h_axi_slave_awready
	wire   [7:0] mm_interconnect_1_hps_0_f2h_axi_slave_awid;     // mm_interconnect_1:hps_0_f2h_axi_slave_awid -> hps_0:f2h_AWID
	wire         mm_interconnect_1_hps_0_f2h_axi_slave_bvalid;   // hps_0:f2h_BVALID -> mm_interconnect_1:hps_0_f2h_axi_slave_bvalid
	wire   [7:0] mm_interconnect_1_hps_0_f2h_axi_slave_wid;      // mm_interconnect_1:hps_0_f2h_axi_slave_wid -> hps_0:f2h_WID
	wire   [1:0] mm_interconnect_1_hps_0_f2h_axi_slave_awlock;   // mm_interconnect_1:hps_0_f2h_axi_slave_awlock -> hps_0:f2h_AWLOCK
	wire   [1:0] mm_interconnect_1_hps_0_f2h_axi_slave_awburst;  // mm_interconnect_1:hps_0_f2h_axi_slave_awburst -> hps_0:f2h_AWBURST
	wire   [1:0] mm_interconnect_1_hps_0_f2h_axi_slave_bresp;    // hps_0:f2h_BRESP -> mm_interconnect_1:hps_0_f2h_axi_slave_bresp
	wire   [4:0] mm_interconnect_1_hps_0_f2h_axi_slave_aruser;   // mm_interconnect_1:hps_0_f2h_axi_slave_aruser -> hps_0:f2h_ARUSER
	wire   [4:0] mm_interconnect_1_hps_0_f2h_axi_slave_awuser;   // mm_interconnect_1:hps_0_f2h_axi_slave_awuser -> hps_0:f2h_AWUSER
	wire   [7:0] mm_interconnect_1_hps_0_f2h_axi_slave_wstrb;    // mm_interconnect_1:hps_0_f2h_axi_slave_wstrb -> hps_0:f2h_WSTRB
	wire         mm_interconnect_1_hps_0_f2h_axi_slave_rvalid;   // hps_0:f2h_RVALID -> mm_interconnect_1:hps_0_f2h_axi_slave_rvalid
	wire   [1:0] mm_interconnect_1_hps_0_f2h_axi_slave_arburst;  // mm_interconnect_1:hps_0_f2h_axi_slave_arburst -> hps_0:f2h_ARBURST
	wire  [63:0] mm_interconnect_1_hps_0_f2h_axi_slave_wdata;    // mm_interconnect_1:hps_0_f2h_axi_slave_wdata -> hps_0:f2h_WDATA
	wire         mm_interconnect_1_hps_0_f2h_axi_slave_wready;   // hps_0:f2h_WREADY -> mm_interconnect_1:hps_0_f2h_axi_slave_wready
	wire  [63:0] mm_interconnect_1_hps_0_f2h_axi_slave_rdata;    // hps_0:f2h_RDATA -> mm_interconnect_1:hps_0_f2h_axi_slave_rdata
	wire  [31:0] mm_interconnect_1_hps_0_f2h_axi_slave_araddr;   // mm_interconnect_1:hps_0_f2h_axi_slave_araddr -> hps_0:f2h_ARADDR
	wire   [3:0] mm_interconnect_1_hps_0_f2h_axi_slave_arcache;  // mm_interconnect_1:hps_0_f2h_axi_slave_arcache -> hps_0:f2h_ARCACHE
	wire   [3:0] mm_interconnect_1_hps_0_f2h_axi_slave_awlen;    // mm_interconnect_1:hps_0_f2h_axi_slave_awlen -> hps_0:f2h_AWLEN
	wire  [31:0] mm_interconnect_1_hps_0_f2h_axi_slave_awaddr;   // mm_interconnect_1:hps_0_f2h_axi_slave_awaddr -> hps_0:f2h_AWADDR
	wire   [7:0] mm_interconnect_1_hps_0_f2h_axi_slave_rid;      // hps_0:f2h_RID -> mm_interconnect_1:hps_0_f2h_axi_slave_rid
	wire         mm_interconnect_1_hps_0_f2h_axi_slave_wvalid;   // mm_interconnect_1:hps_0_f2h_axi_slave_wvalid -> hps_0:f2h_WVALID
	wire   [1:0] mm_interconnect_1_hps_0_f2h_axi_slave_rresp;    // hps_0:f2h_RRESP -> mm_interconnect_1:hps_0_f2h_axi_slave_rresp
	wire         mm_interconnect_1_hps_0_f2h_axi_slave_wlast;    // mm_interconnect_1:hps_0_f2h_axi_slave_wlast -> hps_0:f2h_WLAST
	wire         mm_interconnect_1_hps_0_f2h_axi_slave_rlast;    // hps_0:f2h_RLAST -> mm_interconnect_1:hps_0_f2h_axi_slave_rlast
	wire         hps_0_h2f_reset_reset;                          // hps_0:h2f_rst_n -> rst_controller:reset_in0

	soc_ethond_hps_0 #(
		.F2S_Width (2),
		.S2F_Width (1)
	) hps_0 (
		.h2f_loan_in               (hps_loan_io_in),                                //    h2f_loan_io.in
		.h2f_loan_out              (hps_loan_io_out),                               //               .out
		.h2f_loan_oe               (hps_loan_io_oe),                                //               .oe
		.mem_a                     (memory_mem_a),                                  //         memory.mem_a
		.mem_ba                    (memory_mem_ba),                                 //               .mem_ba
		.mem_ck                    (memory_mem_ck),                                 //               .mem_ck
		.mem_ck_n                  (memory_mem_ck_n),                               //               .mem_ck_n
		.mem_cke                   (memory_mem_cke),                                //               .mem_cke
		.mem_cs_n                  (memory_mem_cs_n),                               //               .mem_cs_n
		.mem_ras_n                 (memory_mem_ras_n),                              //               .mem_ras_n
		.mem_cas_n                 (memory_mem_cas_n),                              //               .mem_cas_n
		.mem_we_n                  (memory_mem_we_n),                               //               .mem_we_n
		.mem_reset_n               (memory_mem_reset_n),                            //               .mem_reset_n
		.mem_dq                    (memory_mem_dq),                                 //               .mem_dq
		.mem_dqs                   (memory_mem_dqs),                                //               .mem_dqs
		.mem_dqs_n                 (memory_mem_dqs_n),                              //               .mem_dqs_n
		.mem_odt                   (memory_mem_odt),                                //               .mem_odt
		.mem_dm                    (memory_mem_dm),                                 //               .mem_dm
		.oct_rzqin                 (memory_oct_rzqin),                              //               .oct_rzqin
		.hps_io_emac1_inst_TX_CLK  (hps_io_hps_io_emac1_inst_TX_CLK),               //         hps_io.hps_io_emac1_inst_TX_CLK
		.hps_io_emac1_inst_TXD0    (hps_io_hps_io_emac1_inst_TXD0),                 //               .hps_io_emac1_inst_TXD0
		.hps_io_emac1_inst_TXD1    (hps_io_hps_io_emac1_inst_TXD1),                 //               .hps_io_emac1_inst_TXD1
		.hps_io_emac1_inst_TXD2    (hps_io_hps_io_emac1_inst_TXD2),                 //               .hps_io_emac1_inst_TXD2
		.hps_io_emac1_inst_TXD3    (hps_io_hps_io_emac1_inst_TXD3),                 //               .hps_io_emac1_inst_TXD3
		.hps_io_emac1_inst_RXD0    (hps_io_hps_io_emac1_inst_RXD0),                 //               .hps_io_emac1_inst_RXD0
		.hps_io_emac1_inst_MDIO    (hps_io_hps_io_emac1_inst_MDIO),                 //               .hps_io_emac1_inst_MDIO
		.hps_io_emac1_inst_MDC     (hps_io_hps_io_emac1_inst_MDC),                  //               .hps_io_emac1_inst_MDC
		.hps_io_emac1_inst_RX_CTL  (hps_io_hps_io_emac1_inst_RX_CTL),               //               .hps_io_emac1_inst_RX_CTL
		.hps_io_emac1_inst_TX_CTL  (hps_io_hps_io_emac1_inst_TX_CTL),               //               .hps_io_emac1_inst_TX_CTL
		.hps_io_emac1_inst_RX_CLK  (hps_io_hps_io_emac1_inst_RX_CLK),               //               .hps_io_emac1_inst_RX_CLK
		.hps_io_emac1_inst_RXD1    (hps_io_hps_io_emac1_inst_RXD1),                 //               .hps_io_emac1_inst_RXD1
		.hps_io_emac1_inst_RXD2    (hps_io_hps_io_emac1_inst_RXD2),                 //               .hps_io_emac1_inst_RXD2
		.hps_io_emac1_inst_RXD3    (hps_io_hps_io_emac1_inst_RXD3),                 //               .hps_io_emac1_inst_RXD3
		.hps_io_qspi_inst_IO0      (hps_io_hps_io_qspi_inst_IO0),                   //               .hps_io_qspi_inst_IO0
		.hps_io_qspi_inst_IO1      (hps_io_hps_io_qspi_inst_IO1),                   //               .hps_io_qspi_inst_IO1
		.hps_io_qspi_inst_IO2      (hps_io_hps_io_qspi_inst_IO2),                   //               .hps_io_qspi_inst_IO2
		.hps_io_qspi_inst_IO3      (hps_io_hps_io_qspi_inst_IO3),                   //               .hps_io_qspi_inst_IO3
		.hps_io_qspi_inst_SS0      (hps_io_hps_io_qspi_inst_SS0),                   //               .hps_io_qspi_inst_SS0
		.hps_io_qspi_inst_CLK      (hps_io_hps_io_qspi_inst_CLK),                   //               .hps_io_qspi_inst_CLK
		.hps_io_sdio_inst_CMD      (hps_io_hps_io_sdio_inst_CMD),                   //               .hps_io_sdio_inst_CMD
		.hps_io_sdio_inst_D0       (hps_io_hps_io_sdio_inst_D0),                    //               .hps_io_sdio_inst_D0
		.hps_io_sdio_inst_D1       (hps_io_hps_io_sdio_inst_D1),                    //               .hps_io_sdio_inst_D1
		.hps_io_sdio_inst_CLK      (hps_io_hps_io_sdio_inst_CLK),                   //               .hps_io_sdio_inst_CLK
		.hps_io_sdio_inst_D2       (hps_io_hps_io_sdio_inst_D2),                    //               .hps_io_sdio_inst_D2
		.hps_io_sdio_inst_D3       (hps_io_hps_io_sdio_inst_D3),                    //               .hps_io_sdio_inst_D3
		.hps_io_usb1_inst_D0       (hps_io_hps_io_usb1_inst_D0),                    //               .hps_io_usb1_inst_D0
		.hps_io_usb1_inst_D1       (hps_io_hps_io_usb1_inst_D1),                    //               .hps_io_usb1_inst_D1
		.hps_io_usb1_inst_D2       (hps_io_hps_io_usb1_inst_D2),                    //               .hps_io_usb1_inst_D2
		.hps_io_usb1_inst_D3       (hps_io_hps_io_usb1_inst_D3),                    //               .hps_io_usb1_inst_D3
		.hps_io_usb1_inst_D4       (hps_io_hps_io_usb1_inst_D4),                    //               .hps_io_usb1_inst_D4
		.hps_io_usb1_inst_D5       (hps_io_hps_io_usb1_inst_D5),                    //               .hps_io_usb1_inst_D5
		.hps_io_usb1_inst_D6       (hps_io_hps_io_usb1_inst_D6),                    //               .hps_io_usb1_inst_D6
		.hps_io_usb1_inst_D7       (hps_io_hps_io_usb1_inst_D7),                    //               .hps_io_usb1_inst_D7
		.hps_io_usb1_inst_CLK      (hps_io_hps_io_usb1_inst_CLK),                   //               .hps_io_usb1_inst_CLK
		.hps_io_usb1_inst_STP      (hps_io_hps_io_usb1_inst_STP),                   //               .hps_io_usb1_inst_STP
		.hps_io_usb1_inst_DIR      (hps_io_hps_io_usb1_inst_DIR),                   //               .hps_io_usb1_inst_DIR
		.hps_io_usb1_inst_NXT      (hps_io_hps_io_usb1_inst_NXT),                   //               .hps_io_usb1_inst_NXT
		.hps_io_uart0_inst_RX      (hps_io_hps_io_uart0_inst_RX),                   //               .hps_io_uart0_inst_RX
		.hps_io_uart0_inst_TX      (hps_io_hps_io_uart0_inst_TX),                   //               .hps_io_uart0_inst_TX
		.hps_io_i2c0_inst_SDA      (hps_io_hps_io_i2c0_inst_SDA),                   //               .hps_io_i2c0_inst_SDA
		.hps_io_i2c0_inst_SCL      (hps_io_hps_io_i2c0_inst_SCL),                   //               .hps_io_i2c0_inst_SCL
		.hps_io_gpio_inst_GPIO09   (hps_io_hps_io_gpio_inst_GPIO09),                //               .hps_io_gpio_inst_GPIO09
		.hps_io_gpio_inst_GPIO37   (hps_io_hps_io_gpio_inst_GPIO37),                //               .hps_io_gpio_inst_GPIO37
		.hps_io_gpio_inst_GPIO44   (hps_io_hps_io_gpio_inst_GPIO44),                //               .hps_io_gpio_inst_GPIO44
		.hps_io_gpio_inst_GPIO48   (hps_io_hps_io_gpio_inst_GPIO48),                //               .hps_io_gpio_inst_GPIO48
		.hps_io_gpio_inst_GPIO52   (hps_io_hps_io_gpio_inst_GPIO52),                //               .hps_io_gpio_inst_GPIO52
		.hps_io_gpio_inst_GPIO65   (hps_io_hps_io_gpio_inst_GPIO65),                //               .hps_io_gpio_inst_GPIO65
		.hps_io_gpio_inst_LOANIO58 (hps_io_hps_io_gpio_inst_LOANIO58),              //               .hps_io_gpio_inst_LOANIO58
		.h2f_rst_n                 (hps_0_h2f_reset_reset),                         //      h2f_reset.reset_n
		.h2f_axi_clk               (sys_clk_clk),                                   //  h2f_axi_clock.clk
		.h2f_AWID                  (hps_0_h2f_axi_master_awid),                     // h2f_axi_master.awid
		.h2f_AWADDR                (hps_0_h2f_axi_master_awaddr),                   //               .awaddr
		.h2f_AWLEN                 (hps_0_h2f_axi_master_awlen),                    //               .awlen
		.h2f_AWSIZE                (hps_0_h2f_axi_master_awsize),                   //               .awsize
		.h2f_AWBURST               (hps_0_h2f_axi_master_awburst),                  //               .awburst
		.h2f_AWLOCK                (hps_0_h2f_axi_master_awlock),                   //               .awlock
		.h2f_AWCACHE               (hps_0_h2f_axi_master_awcache),                  //               .awcache
		.h2f_AWPROT                (hps_0_h2f_axi_master_awprot),                   //               .awprot
		.h2f_AWVALID               (hps_0_h2f_axi_master_awvalid),                  //               .awvalid
		.h2f_AWREADY               (hps_0_h2f_axi_master_awready),                  //               .awready
		.h2f_WID                   (hps_0_h2f_axi_master_wid),                      //               .wid
		.h2f_WDATA                 (hps_0_h2f_axi_master_wdata),                    //               .wdata
		.h2f_WSTRB                 (hps_0_h2f_axi_master_wstrb),                    //               .wstrb
		.h2f_WLAST                 (hps_0_h2f_axi_master_wlast),                    //               .wlast
		.h2f_WVALID                (hps_0_h2f_axi_master_wvalid),                   //               .wvalid
		.h2f_WREADY                (hps_0_h2f_axi_master_wready),                   //               .wready
		.h2f_BID                   (hps_0_h2f_axi_master_bid),                      //               .bid
		.h2f_BRESP                 (hps_0_h2f_axi_master_bresp),                    //               .bresp
		.h2f_BVALID                (hps_0_h2f_axi_master_bvalid),                   //               .bvalid
		.h2f_BREADY                (hps_0_h2f_axi_master_bready),                   //               .bready
		.h2f_ARID                  (hps_0_h2f_axi_master_arid),                     //               .arid
		.h2f_ARADDR                (hps_0_h2f_axi_master_araddr),                   //               .araddr
		.h2f_ARLEN                 (hps_0_h2f_axi_master_arlen),                    //               .arlen
		.h2f_ARSIZE                (hps_0_h2f_axi_master_arsize),                   //               .arsize
		.h2f_ARBURST               (hps_0_h2f_axi_master_arburst),                  //               .arburst
		.h2f_ARLOCK                (hps_0_h2f_axi_master_arlock),                   //               .arlock
		.h2f_ARCACHE               (hps_0_h2f_axi_master_arcache),                  //               .arcache
		.h2f_ARPROT                (hps_0_h2f_axi_master_arprot),                   //               .arprot
		.h2f_ARVALID               (hps_0_h2f_axi_master_arvalid),                  //               .arvalid
		.h2f_ARREADY               (hps_0_h2f_axi_master_arready),                  //               .arready
		.h2f_RID                   (hps_0_h2f_axi_master_rid),                      //               .rid
		.h2f_RDATA                 (hps_0_h2f_axi_master_rdata),                    //               .rdata
		.h2f_RRESP                 (hps_0_h2f_axi_master_rresp),                    //               .rresp
		.h2f_RLAST                 (hps_0_h2f_axi_master_rlast),                    //               .rlast
		.h2f_RVALID                (hps_0_h2f_axi_master_rvalid),                   //               .rvalid
		.h2f_RREADY                (hps_0_h2f_axi_master_rready),                   //               .rready
		.f2h_axi_clk               (sys_clk_clk),                                   //  f2h_axi_clock.clk
		.f2h_AWID                  (mm_interconnect_1_hps_0_f2h_axi_slave_awid),    //  f2h_axi_slave.awid
		.f2h_AWADDR                (mm_interconnect_1_hps_0_f2h_axi_slave_awaddr),  //               .awaddr
		.f2h_AWLEN                 (mm_interconnect_1_hps_0_f2h_axi_slave_awlen),   //               .awlen
		.f2h_AWSIZE                (mm_interconnect_1_hps_0_f2h_axi_slave_awsize),  //               .awsize
		.f2h_AWBURST               (mm_interconnect_1_hps_0_f2h_axi_slave_awburst), //               .awburst
		.f2h_AWLOCK                (mm_interconnect_1_hps_0_f2h_axi_slave_awlock),  //               .awlock
		.f2h_AWCACHE               (mm_interconnect_1_hps_0_f2h_axi_slave_awcache), //               .awcache
		.f2h_AWPROT                (mm_interconnect_1_hps_0_f2h_axi_slave_awprot),  //               .awprot
		.f2h_AWVALID               (mm_interconnect_1_hps_0_f2h_axi_slave_awvalid), //               .awvalid
		.f2h_AWREADY               (mm_interconnect_1_hps_0_f2h_axi_slave_awready), //               .awready
		.f2h_AWUSER                (mm_interconnect_1_hps_0_f2h_axi_slave_awuser),  //               .awuser
		.f2h_WID                   (mm_interconnect_1_hps_0_f2h_axi_slave_wid),     //               .wid
		.f2h_WDATA                 (mm_interconnect_1_hps_0_f2h_axi_slave_wdata),   //               .wdata
		.f2h_WSTRB                 (mm_interconnect_1_hps_0_f2h_axi_slave_wstrb),   //               .wstrb
		.f2h_WLAST                 (mm_interconnect_1_hps_0_f2h_axi_slave_wlast),   //               .wlast
		.f2h_WVALID                (mm_interconnect_1_hps_0_f2h_axi_slave_wvalid),  //               .wvalid
		.f2h_WREADY                (mm_interconnect_1_hps_0_f2h_axi_slave_wready),  //               .wready
		.f2h_BID                   (mm_interconnect_1_hps_0_f2h_axi_slave_bid),     //               .bid
		.f2h_BRESP                 (mm_interconnect_1_hps_0_f2h_axi_slave_bresp),   //               .bresp
		.f2h_BVALID                (mm_interconnect_1_hps_0_f2h_axi_slave_bvalid),  //               .bvalid
		.f2h_BREADY                (mm_interconnect_1_hps_0_f2h_axi_slave_bready),  //               .bready
		.f2h_ARID                  (mm_interconnect_1_hps_0_f2h_axi_slave_arid),    //               .arid
		.f2h_ARADDR                (mm_interconnect_1_hps_0_f2h_axi_slave_araddr),  //               .araddr
		.f2h_ARLEN                 (mm_interconnect_1_hps_0_f2h_axi_slave_arlen),   //               .arlen
		.f2h_ARSIZE                (mm_interconnect_1_hps_0_f2h_axi_slave_arsize),  //               .arsize
		.f2h_ARBURST               (mm_interconnect_1_hps_0_f2h_axi_slave_arburst), //               .arburst
		.f2h_ARLOCK                (mm_interconnect_1_hps_0_f2h_axi_slave_arlock),  //               .arlock
		.f2h_ARCACHE               (mm_interconnect_1_hps_0_f2h_axi_slave_arcache), //               .arcache
		.f2h_ARPROT                (mm_interconnect_1_hps_0_f2h_axi_slave_arprot),  //               .arprot
		.f2h_ARVALID               (mm_interconnect_1_hps_0_f2h_axi_slave_arvalid), //               .arvalid
		.f2h_ARREADY               (mm_interconnect_1_hps_0_f2h_axi_slave_arready), //               .arready
		.f2h_ARUSER                (mm_interconnect_1_hps_0_f2h_axi_slave_aruser),  //               .aruser
		.f2h_RID                   (mm_interconnect_1_hps_0_f2h_axi_slave_rid),     //               .rid
		.f2h_RDATA                 (mm_interconnect_1_hps_0_f2h_axi_slave_rdata),   //               .rdata
		.f2h_RRESP                 (mm_interconnect_1_hps_0_f2h_axi_slave_rresp),   //               .rresp
		.f2h_RLAST                 (mm_interconnect_1_hps_0_f2h_axi_slave_rlast),   //               .rlast
		.f2h_RVALID                (mm_interconnect_1_hps_0_f2h_axi_slave_rvalid),  //               .rvalid
		.f2h_RREADY                (mm_interconnect_1_hps_0_f2h_axi_slave_rready),  //               .rready
		.f2h_irq_p0                (irq0_irq),                                      //       f2h_irq0.irq
		.f2h_irq_p1                (irq1_irq)                                       //       f2h_irq1.irq
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (32),
		.SYMBOL_WIDTH      (8),
		.HDL_ADDR_WIDTH    (13),
		.BURSTCOUNT_WIDTH  (1),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) mm_bridge_0 (
		.clk              (sys_clk_clk),                                    //   clk.clk
		.reset            (sys_rst_reset),                                  // reset.reset
		.s0_waitrequest   (mm_interconnect_0_mm_bridge_0_s0_waitrequest),   //    s0.waitrequest
		.s0_readdata      (mm_interconnect_0_mm_bridge_0_s0_readdata),      //      .readdata
		.s0_readdatavalid (mm_interconnect_0_mm_bridge_0_s0_readdatavalid), //      .readdatavalid
		.s0_burstcount    (mm_interconnect_0_mm_bridge_0_s0_burstcount),    //      .burstcount
		.s0_writedata     (mm_interconnect_0_mm_bridge_0_s0_writedata),     //      .writedata
		.s0_address       (mm_interconnect_0_mm_bridge_0_s0_address),       //      .address
		.s0_write         (mm_interconnect_0_mm_bridge_0_s0_write),         //      .write
		.s0_read          (mm_interconnect_0_mm_bridge_0_s0_read),          //      .read
		.s0_byteenable    (mm_interconnect_0_mm_bridge_0_s0_byteenable),    //      .byteenable
		.s0_debugaccess   (mm_interconnect_0_mm_bridge_0_s0_debugaccess),   //      .debugaccess
		.m0_waitrequest   (csr_waitrequest),                                //    m0.waitrequest
		.m0_readdata      (csr_readdata),                                   //      .readdata
		.m0_readdatavalid (csr_readdatavalid),                              //      .readdatavalid
		.m0_burstcount    (csr_burstcount),                                 //      .burstcount
		.m0_writedata     (csr_writedata),                                  //      .writedata
		.m0_address       (csr_address),                                    //      .address
		.m0_write         (csr_write),                                      //      .write
		.m0_read          (csr_read),                                       //      .read
		.m0_byteenable    (csr_byteenable),                                 //      .byteenable
		.m0_debugaccess   (csr_debugaccess)                                 //      .debugaccess
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (32),
		.SYMBOL_WIDTH      (8),
		.HDL_ADDR_WIDTH    (13),
		.BURSTCOUNT_WIDTH  (1),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) mm_bridge_5 (
		.clk              (sys_clk_clk),                                    //   clk.clk
		.reset            (sys_rst_reset),                                  // reset.reset
		.s0_waitrequest   (mm_interconnect_0_mm_bridge_5_s0_waitrequest),   //    s0.waitrequest
		.s0_readdata      (mm_interconnect_0_mm_bridge_5_s0_readdata),      //      .readdata
		.s0_readdatavalid (mm_interconnect_0_mm_bridge_5_s0_readdatavalid), //      .readdatavalid
		.s0_burstcount    (mm_interconnect_0_mm_bridge_5_s0_burstcount),    //      .burstcount
		.s0_writedata     (mm_interconnect_0_mm_bridge_5_s0_writedata),     //      .writedata
		.s0_address       (mm_interconnect_0_mm_bridge_5_s0_address),       //      .address
		.s0_write         (mm_interconnect_0_mm_bridge_5_s0_write),         //      .write
		.s0_read          (mm_interconnect_0_mm_bridge_5_s0_read),          //      .read
		.s0_byteenable    (mm_interconnect_0_mm_bridge_5_s0_byteenable),    //      .byteenable
		.s0_debugaccess   (mm_interconnect_0_mm_bridge_5_s0_debugaccess),   //      .debugaccess
		.m0_waitrequest   (netdma_csr0_waitrequest),                        //    m0.waitrequest
		.m0_readdata      (netdma_csr0_readdata),                           //      .readdata
		.m0_readdatavalid (netdma_csr0_readdatavalid),                      //      .readdatavalid
		.m0_burstcount    (netdma_csr0_burstcount),                         //      .burstcount
		.m0_writedata     (netdma_csr0_writedata),                          //      .writedata
		.m0_address       (netdma_csr0_address),                            //      .address
		.m0_write         (netdma_csr0_write),                              //      .write
		.m0_read          (netdma_csr0_read),                               //      .read
		.m0_byteenable    (netdma_csr0_byteenable),                         //      .byteenable
		.m0_debugaccess   (netdma_csr0_debugaccess)                         //      .debugaccess
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (32),
		.SYMBOL_WIDTH      (8),
		.HDL_ADDR_WIDTH    (13),
		.BURSTCOUNT_WIDTH  (1),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) mm_bridge_6 (
		.clk              (sys_clk_clk),                                    //   clk.clk
		.reset            (sys_rst_reset),                                  // reset.reset
		.s0_waitrequest   (mm_interconnect_0_mm_bridge_6_s0_waitrequest),   //    s0.waitrequest
		.s0_readdata      (mm_interconnect_0_mm_bridge_6_s0_readdata),      //      .readdata
		.s0_readdatavalid (mm_interconnect_0_mm_bridge_6_s0_readdatavalid), //      .readdatavalid
		.s0_burstcount    (mm_interconnect_0_mm_bridge_6_s0_burstcount),    //      .burstcount
		.s0_writedata     (mm_interconnect_0_mm_bridge_6_s0_writedata),     //      .writedata
		.s0_address       (mm_interconnect_0_mm_bridge_6_s0_address),       //      .address
		.s0_write         (mm_interconnect_0_mm_bridge_6_s0_write),         //      .write
		.s0_read          (mm_interconnect_0_mm_bridge_6_s0_read),          //      .read
		.s0_byteenable    (mm_interconnect_0_mm_bridge_6_s0_byteenable),    //      .byteenable
		.s0_debugaccess   (mm_interconnect_0_mm_bridge_6_s0_debugaccess),   //      .debugaccess
		.m0_waitrequest   (netdma_csr1_waitrequest),                        //    m0.waitrequest
		.m0_readdata      (netdma_csr1_readdata),                           //      .readdata
		.m0_readdatavalid (netdma_csr1_readdatavalid),                      //      .readdatavalid
		.m0_burstcount    (netdma_csr1_burstcount),                         //      .burstcount
		.m0_writedata     (netdma_csr1_writedata),                          //      .writedata
		.m0_address       (netdma_csr1_address),                            //      .address
		.m0_write         (netdma_csr1_write),                              //      .write
		.m0_read          (netdma_csr1_read),                               //      .read
		.m0_byteenable    (netdma_csr1_byteenable),                         //      .byteenable
		.m0_debugaccess   (netdma_csr1_debugaccess)                         //      .debugaccess
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (64),
		.SYMBOL_WIDTH      (8),
		.HDL_ADDR_WIDTH    (32),
		.BURSTCOUNT_WIDTH  (1),
		.PIPELINE_COMMAND  (0),
		.PIPELINE_RESPONSE (0)
	) mm_bridge_1 (
		.clk              (sys_clk_clk),                  //   clk.clk
		.reset            (sys_rst_reset),                // reset.reset
		.s0_waitrequest   (netdma_read0_waitrequest),     //    s0.waitrequest
		.s0_readdata      (netdma_read0_readdata),        //      .readdata
		.s0_readdatavalid (netdma_read0_readdatavalid),   //      .readdatavalid
		.s0_burstcount    (netdma_read0_burstcount),      //      .burstcount
		.s0_writedata     (netdma_read0_writedata),       //      .writedata
		.s0_address       (netdma_read0_address),         //      .address
		.s0_write         (netdma_read0_write),           //      .write
		.s0_read          (netdma_read0_read),            //      .read
		.s0_byteenable    (netdma_read0_byteenable),      //      .byteenable
		.s0_debugaccess   (netdma_read0_debugaccess),     //      .debugaccess
		.m0_waitrequest   (mm_bridge_1_m0_waitrequest),   //    m0.waitrequest
		.m0_readdata      (mm_bridge_1_m0_readdata),      //      .readdata
		.m0_readdatavalid (mm_bridge_1_m0_readdatavalid), //      .readdatavalid
		.m0_burstcount    (mm_bridge_1_m0_burstcount),    //      .burstcount
		.m0_writedata     (mm_bridge_1_m0_writedata),     //      .writedata
		.m0_address       (mm_bridge_1_m0_address),       //      .address
		.m0_write         (mm_bridge_1_m0_write),         //      .write
		.m0_read          (mm_bridge_1_m0_read),          //      .read
		.m0_byteenable    (mm_bridge_1_m0_byteenable),    //      .byteenable
		.m0_debugaccess   (mm_bridge_1_m0_debugaccess)    //      .debugaccess
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (64),
		.SYMBOL_WIDTH      (8),
		.HDL_ADDR_WIDTH    (32),
		.BURSTCOUNT_WIDTH  (1),
		.PIPELINE_COMMAND  (0),
		.PIPELINE_RESPONSE (0)
	) mm_bridge_2 (
		.clk              (sys_clk_clk),                  //   clk.clk
		.reset            (sys_rst_reset),                // reset.reset
		.s0_waitrequest   (netdma_read1_waitrequest),     //    s0.waitrequest
		.s0_readdata      (netdma_read1_readdata),        //      .readdata
		.s0_readdatavalid (netdma_read1_readdatavalid),   //      .readdatavalid
		.s0_burstcount    (netdma_read1_burstcount),      //      .burstcount
		.s0_writedata     (netdma_read1_writedata),       //      .writedata
		.s0_address       (netdma_read1_address),         //      .address
		.s0_write         (netdma_read1_write),           //      .write
		.s0_read          (netdma_read1_read),            //      .read
		.s0_byteenable    (netdma_read1_byteenable),      //      .byteenable
		.s0_debugaccess   (netdma_read1_debugaccess),     //      .debugaccess
		.m0_waitrequest   (mm_bridge_2_m0_waitrequest),   //    m0.waitrequest
		.m0_readdata      (mm_bridge_2_m0_readdata),      //      .readdata
		.m0_readdatavalid (mm_bridge_2_m0_readdatavalid), //      .readdatavalid
		.m0_burstcount    (mm_bridge_2_m0_burstcount),    //      .burstcount
		.m0_writedata     (mm_bridge_2_m0_writedata),     //      .writedata
		.m0_address       (mm_bridge_2_m0_address),       //      .address
		.m0_write         (mm_bridge_2_m0_write),         //      .write
		.m0_read          (mm_bridge_2_m0_read),          //      .read
		.m0_byteenable    (mm_bridge_2_m0_byteenable),    //      .byteenable
		.m0_debugaccess   (mm_bridge_2_m0_debugaccess)    //      .debugaccess
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (64),
		.SYMBOL_WIDTH      (8),
		.HDL_ADDR_WIDTH    (32),
		.BURSTCOUNT_WIDTH  (1),
		.PIPELINE_COMMAND  (0),
		.PIPELINE_RESPONSE (0)
	) mm_bridge_3 (
		.clk              (sys_clk_clk),                  //   clk.clk
		.reset            (sys_rst_reset),                // reset.reset
		.s0_waitrequest   (netdma_write0_waitrequest),    //    s0.waitrequest
		.s0_readdata      (netdma_write0_readdata),       //      .readdata
		.s0_readdatavalid (netdma_write0_readdatavalid),  //      .readdatavalid
		.s0_burstcount    (netdma_write0_burstcount),     //      .burstcount
		.s0_writedata     (netdma_write0_writedata),      //      .writedata
		.s0_address       (netdma_write0_address),        //      .address
		.s0_write         (netdma_write0_write),          //      .write
		.s0_read          (netdma_write0_read),           //      .read
		.s0_byteenable    (netdma_write0_byteenable),     //      .byteenable
		.s0_debugaccess   (netdma_write0_debugaccess),    //      .debugaccess
		.m0_waitrequest   (mm_bridge_3_m0_waitrequest),   //    m0.waitrequest
		.m0_readdata      (mm_bridge_3_m0_readdata),      //      .readdata
		.m0_readdatavalid (mm_bridge_3_m0_readdatavalid), //      .readdatavalid
		.m0_burstcount    (mm_bridge_3_m0_burstcount),    //      .burstcount
		.m0_writedata     (mm_bridge_3_m0_writedata),     //      .writedata
		.m0_address       (mm_bridge_3_m0_address),       //      .address
		.m0_write         (mm_bridge_3_m0_write),         //      .write
		.m0_read          (mm_bridge_3_m0_read),          //      .read
		.m0_byteenable    (mm_bridge_3_m0_byteenable),    //      .byteenable
		.m0_debugaccess   (mm_bridge_3_m0_debugaccess)    //      .debugaccess
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (64),
		.SYMBOL_WIDTH      (8),
		.HDL_ADDR_WIDTH    (32),
		.BURSTCOUNT_WIDTH  (1),
		.PIPELINE_COMMAND  (0),
		.PIPELINE_RESPONSE (0)
	) mm_bridge_4 (
		.clk              (sys_clk_clk),                  //   clk.clk
		.reset            (sys_rst_reset),                // reset.reset
		.s0_waitrequest   (netdma_write1_waitrequest),    //    s0.waitrequest
		.s0_readdata      (netdma_write1_readdata),       //      .readdata
		.s0_readdatavalid (netdma_write1_readdatavalid),  //      .readdatavalid
		.s0_burstcount    (netdma_write1_burstcount),     //      .burstcount
		.s0_writedata     (netdma_write1_writedata),      //      .writedata
		.s0_address       (netdma_write1_address),        //      .address
		.s0_write         (netdma_write1_write),          //      .write
		.s0_read          (netdma_write1_read),           //      .read
		.s0_byteenable    (netdma_write1_byteenable),     //      .byteenable
		.s0_debugaccess   (netdma_write1_debugaccess),    //      .debugaccess
		.m0_waitrequest   (mm_bridge_4_m0_waitrequest),   //    m0.waitrequest
		.m0_readdata      (mm_bridge_4_m0_readdata),      //      .readdata
		.m0_readdatavalid (mm_bridge_4_m0_readdatavalid), //      .readdatavalid
		.m0_burstcount    (mm_bridge_4_m0_burstcount),    //      .burstcount
		.m0_writedata     (mm_bridge_4_m0_writedata),     //      .writedata
		.m0_address       (mm_bridge_4_m0_address),       //      .address
		.m0_write         (mm_bridge_4_m0_write),         //      .write
		.m0_read          (mm_bridge_4_m0_read),          //      .read
		.m0_byteenable    (mm_bridge_4_m0_byteenable),    //      .byteenable
		.m0_debugaccess   (mm_bridge_4_m0_debugaccess)    //      .debugaccess
	);

	soc_ethond_mm_interconnect_0 mm_interconnect_0 (
		.hps_0_h2f_axi_master_awid                     (hps_0_h2f_axi_master_awid),                      //                    hps_0_h2f_axi_master.awid
		.hps_0_h2f_axi_master_awaddr                   (hps_0_h2f_axi_master_awaddr),                    //                                        .awaddr
		.hps_0_h2f_axi_master_awlen                    (hps_0_h2f_axi_master_awlen),                     //                                        .awlen
		.hps_0_h2f_axi_master_awsize                   (hps_0_h2f_axi_master_awsize),                    //                                        .awsize
		.hps_0_h2f_axi_master_awburst                  (hps_0_h2f_axi_master_awburst),                   //                                        .awburst
		.hps_0_h2f_axi_master_awlock                   (hps_0_h2f_axi_master_awlock),                    //                                        .awlock
		.hps_0_h2f_axi_master_awcache                  (hps_0_h2f_axi_master_awcache),                   //                                        .awcache
		.hps_0_h2f_axi_master_awprot                   (hps_0_h2f_axi_master_awprot),                    //                                        .awprot
		.hps_0_h2f_axi_master_awvalid                  (hps_0_h2f_axi_master_awvalid),                   //                                        .awvalid
		.hps_0_h2f_axi_master_awready                  (hps_0_h2f_axi_master_awready),                   //                                        .awready
		.hps_0_h2f_axi_master_wid                      (hps_0_h2f_axi_master_wid),                       //                                        .wid
		.hps_0_h2f_axi_master_wdata                    (hps_0_h2f_axi_master_wdata),                     //                                        .wdata
		.hps_0_h2f_axi_master_wstrb                    (hps_0_h2f_axi_master_wstrb),                     //                                        .wstrb
		.hps_0_h2f_axi_master_wlast                    (hps_0_h2f_axi_master_wlast),                     //                                        .wlast
		.hps_0_h2f_axi_master_wvalid                   (hps_0_h2f_axi_master_wvalid),                    //                                        .wvalid
		.hps_0_h2f_axi_master_wready                   (hps_0_h2f_axi_master_wready),                    //                                        .wready
		.hps_0_h2f_axi_master_bid                      (hps_0_h2f_axi_master_bid),                       //                                        .bid
		.hps_0_h2f_axi_master_bresp                    (hps_0_h2f_axi_master_bresp),                     //                                        .bresp
		.hps_0_h2f_axi_master_bvalid                   (hps_0_h2f_axi_master_bvalid),                    //                                        .bvalid
		.hps_0_h2f_axi_master_bready                   (hps_0_h2f_axi_master_bready),                    //                                        .bready
		.hps_0_h2f_axi_master_arid                     (hps_0_h2f_axi_master_arid),                      //                                        .arid
		.hps_0_h2f_axi_master_araddr                   (hps_0_h2f_axi_master_araddr),                    //                                        .araddr
		.hps_0_h2f_axi_master_arlen                    (hps_0_h2f_axi_master_arlen),                     //                                        .arlen
		.hps_0_h2f_axi_master_arsize                   (hps_0_h2f_axi_master_arsize),                    //                                        .arsize
		.hps_0_h2f_axi_master_arburst                  (hps_0_h2f_axi_master_arburst),                   //                                        .arburst
		.hps_0_h2f_axi_master_arlock                   (hps_0_h2f_axi_master_arlock),                    //                                        .arlock
		.hps_0_h2f_axi_master_arcache                  (hps_0_h2f_axi_master_arcache),                   //                                        .arcache
		.hps_0_h2f_axi_master_arprot                   (hps_0_h2f_axi_master_arprot),                    //                                        .arprot
		.hps_0_h2f_axi_master_arvalid                  (hps_0_h2f_axi_master_arvalid),                   //                                        .arvalid
		.hps_0_h2f_axi_master_arready                  (hps_0_h2f_axi_master_arready),                   //                                        .arready
		.hps_0_h2f_axi_master_rid                      (hps_0_h2f_axi_master_rid),                       //                                        .rid
		.hps_0_h2f_axi_master_rdata                    (hps_0_h2f_axi_master_rdata),                     //                                        .rdata
		.hps_0_h2f_axi_master_rresp                    (hps_0_h2f_axi_master_rresp),                     //                                        .rresp
		.hps_0_h2f_axi_master_rlast                    (hps_0_h2f_axi_master_rlast),                     //                                        .rlast
		.hps_0_h2f_axi_master_rvalid                   (hps_0_h2f_axi_master_rvalid),                    //                                        .rvalid
		.hps_0_h2f_axi_master_rready                   (hps_0_h2f_axi_master_rready),                    //                                        .rready
		.clock_bridge_0_out_clk_clk                    (sys_clk_clk),                                    //                  clock_bridge_0_out_clk.clk
		.mm_bridge_5_reset_reset_bridge_in_reset_reset (sys_rst_reset),                                  // mm_bridge_5_reset_reset_bridge_in_reset.reset
		.mm_bridge_0_s0_address                        (mm_interconnect_0_mm_bridge_0_s0_address),       //                          mm_bridge_0_s0.address
		.mm_bridge_0_s0_write                          (mm_interconnect_0_mm_bridge_0_s0_write),         //                                        .write
		.mm_bridge_0_s0_read                           (mm_interconnect_0_mm_bridge_0_s0_read),          //                                        .read
		.mm_bridge_0_s0_readdata                       (mm_interconnect_0_mm_bridge_0_s0_readdata),      //                                        .readdata
		.mm_bridge_0_s0_writedata                      (mm_interconnect_0_mm_bridge_0_s0_writedata),     //                                        .writedata
		.mm_bridge_0_s0_burstcount                     (mm_interconnect_0_mm_bridge_0_s0_burstcount),    //                                        .burstcount
		.mm_bridge_0_s0_byteenable                     (mm_interconnect_0_mm_bridge_0_s0_byteenable),    //                                        .byteenable
		.mm_bridge_0_s0_readdatavalid                  (mm_interconnect_0_mm_bridge_0_s0_readdatavalid), //                                        .readdatavalid
		.mm_bridge_0_s0_waitrequest                    (mm_interconnect_0_mm_bridge_0_s0_waitrequest),   //                                        .waitrequest
		.mm_bridge_0_s0_debugaccess                    (mm_interconnect_0_mm_bridge_0_s0_debugaccess),   //                                        .debugaccess
		.mm_bridge_5_s0_address                        (mm_interconnect_0_mm_bridge_5_s0_address),       //                          mm_bridge_5_s0.address
		.mm_bridge_5_s0_write                          (mm_interconnect_0_mm_bridge_5_s0_write),         //                                        .write
		.mm_bridge_5_s0_read                           (mm_interconnect_0_mm_bridge_5_s0_read),          //                                        .read
		.mm_bridge_5_s0_readdata                       (mm_interconnect_0_mm_bridge_5_s0_readdata),      //                                        .readdata
		.mm_bridge_5_s0_writedata                      (mm_interconnect_0_mm_bridge_5_s0_writedata),     //                                        .writedata
		.mm_bridge_5_s0_burstcount                     (mm_interconnect_0_mm_bridge_5_s0_burstcount),    //                                        .burstcount
		.mm_bridge_5_s0_byteenable                     (mm_interconnect_0_mm_bridge_5_s0_byteenable),    //                                        .byteenable
		.mm_bridge_5_s0_readdatavalid                  (mm_interconnect_0_mm_bridge_5_s0_readdatavalid), //                                        .readdatavalid
		.mm_bridge_5_s0_waitrequest                    (mm_interconnect_0_mm_bridge_5_s0_waitrequest),   //                                        .waitrequest
		.mm_bridge_5_s0_debugaccess                    (mm_interconnect_0_mm_bridge_5_s0_debugaccess),   //                                        .debugaccess
		.mm_bridge_6_s0_address                        (mm_interconnect_0_mm_bridge_6_s0_address),       //                          mm_bridge_6_s0.address
		.mm_bridge_6_s0_write                          (mm_interconnect_0_mm_bridge_6_s0_write),         //                                        .write
		.mm_bridge_6_s0_read                           (mm_interconnect_0_mm_bridge_6_s0_read),          //                                        .read
		.mm_bridge_6_s0_readdata                       (mm_interconnect_0_mm_bridge_6_s0_readdata),      //                                        .readdata
		.mm_bridge_6_s0_writedata                      (mm_interconnect_0_mm_bridge_6_s0_writedata),     //                                        .writedata
		.mm_bridge_6_s0_burstcount                     (mm_interconnect_0_mm_bridge_6_s0_burstcount),    //                                        .burstcount
		.mm_bridge_6_s0_byteenable                     (mm_interconnect_0_mm_bridge_6_s0_byteenable),    //                                        .byteenable
		.mm_bridge_6_s0_readdatavalid                  (mm_interconnect_0_mm_bridge_6_s0_readdatavalid), //                                        .readdatavalid
		.mm_bridge_6_s0_waitrequest                    (mm_interconnect_0_mm_bridge_6_s0_waitrequest),   //                                        .waitrequest
		.mm_bridge_6_s0_debugaccess                    (mm_interconnect_0_mm_bridge_6_s0_debugaccess)    //                                        .debugaccess
	);

	soc_ethond_mm_interconnect_1 mm_interconnect_1 (
		.hps_0_f2h_axi_slave_awid                      (mm_interconnect_1_hps_0_f2h_axi_slave_awid),    //                     hps_0_f2h_axi_slave.awid
		.hps_0_f2h_axi_slave_awaddr                    (mm_interconnect_1_hps_0_f2h_axi_slave_awaddr),  //                                        .awaddr
		.hps_0_f2h_axi_slave_awlen                     (mm_interconnect_1_hps_0_f2h_axi_slave_awlen),   //                                        .awlen
		.hps_0_f2h_axi_slave_awsize                    (mm_interconnect_1_hps_0_f2h_axi_slave_awsize),  //                                        .awsize
		.hps_0_f2h_axi_slave_awburst                   (mm_interconnect_1_hps_0_f2h_axi_slave_awburst), //                                        .awburst
		.hps_0_f2h_axi_slave_awlock                    (mm_interconnect_1_hps_0_f2h_axi_slave_awlock),  //                                        .awlock
		.hps_0_f2h_axi_slave_awcache                   (mm_interconnect_1_hps_0_f2h_axi_slave_awcache), //                                        .awcache
		.hps_0_f2h_axi_slave_awprot                    (mm_interconnect_1_hps_0_f2h_axi_slave_awprot),  //                                        .awprot
		.hps_0_f2h_axi_slave_awuser                    (mm_interconnect_1_hps_0_f2h_axi_slave_awuser),  //                                        .awuser
		.hps_0_f2h_axi_slave_awvalid                   (mm_interconnect_1_hps_0_f2h_axi_slave_awvalid), //                                        .awvalid
		.hps_0_f2h_axi_slave_awready                   (mm_interconnect_1_hps_0_f2h_axi_slave_awready), //                                        .awready
		.hps_0_f2h_axi_slave_wid                       (mm_interconnect_1_hps_0_f2h_axi_slave_wid),     //                                        .wid
		.hps_0_f2h_axi_slave_wdata                     (mm_interconnect_1_hps_0_f2h_axi_slave_wdata),   //                                        .wdata
		.hps_0_f2h_axi_slave_wstrb                     (mm_interconnect_1_hps_0_f2h_axi_slave_wstrb),   //                                        .wstrb
		.hps_0_f2h_axi_slave_wlast                     (mm_interconnect_1_hps_0_f2h_axi_slave_wlast),   //                                        .wlast
		.hps_0_f2h_axi_slave_wvalid                    (mm_interconnect_1_hps_0_f2h_axi_slave_wvalid),  //                                        .wvalid
		.hps_0_f2h_axi_slave_wready                    (mm_interconnect_1_hps_0_f2h_axi_slave_wready),  //                                        .wready
		.hps_0_f2h_axi_slave_bid                       (mm_interconnect_1_hps_0_f2h_axi_slave_bid),     //                                        .bid
		.hps_0_f2h_axi_slave_bresp                     (mm_interconnect_1_hps_0_f2h_axi_slave_bresp),   //                                        .bresp
		.hps_0_f2h_axi_slave_bvalid                    (mm_interconnect_1_hps_0_f2h_axi_slave_bvalid),  //                                        .bvalid
		.hps_0_f2h_axi_slave_bready                    (mm_interconnect_1_hps_0_f2h_axi_slave_bready),  //                                        .bready
		.hps_0_f2h_axi_slave_arid                      (mm_interconnect_1_hps_0_f2h_axi_slave_arid),    //                                        .arid
		.hps_0_f2h_axi_slave_araddr                    (mm_interconnect_1_hps_0_f2h_axi_slave_araddr),  //                                        .araddr
		.hps_0_f2h_axi_slave_arlen                     (mm_interconnect_1_hps_0_f2h_axi_slave_arlen),   //                                        .arlen
		.hps_0_f2h_axi_slave_arsize                    (mm_interconnect_1_hps_0_f2h_axi_slave_arsize),  //                                        .arsize
		.hps_0_f2h_axi_slave_arburst                   (mm_interconnect_1_hps_0_f2h_axi_slave_arburst), //                                        .arburst
		.hps_0_f2h_axi_slave_arlock                    (mm_interconnect_1_hps_0_f2h_axi_slave_arlock),  //                                        .arlock
		.hps_0_f2h_axi_slave_arcache                   (mm_interconnect_1_hps_0_f2h_axi_slave_arcache), //                                        .arcache
		.hps_0_f2h_axi_slave_arprot                    (mm_interconnect_1_hps_0_f2h_axi_slave_arprot),  //                                        .arprot
		.hps_0_f2h_axi_slave_aruser                    (mm_interconnect_1_hps_0_f2h_axi_slave_aruser),  //                                        .aruser
		.hps_0_f2h_axi_slave_arvalid                   (mm_interconnect_1_hps_0_f2h_axi_slave_arvalid), //                                        .arvalid
		.hps_0_f2h_axi_slave_arready                   (mm_interconnect_1_hps_0_f2h_axi_slave_arready), //                                        .arready
		.hps_0_f2h_axi_slave_rid                       (mm_interconnect_1_hps_0_f2h_axi_slave_rid),     //                                        .rid
		.hps_0_f2h_axi_slave_rdata                     (mm_interconnect_1_hps_0_f2h_axi_slave_rdata),   //                                        .rdata
		.hps_0_f2h_axi_slave_rresp                     (mm_interconnect_1_hps_0_f2h_axi_slave_rresp),   //                                        .rresp
		.hps_0_f2h_axi_slave_rlast                     (mm_interconnect_1_hps_0_f2h_axi_slave_rlast),   //                                        .rlast
		.hps_0_f2h_axi_slave_rvalid                    (mm_interconnect_1_hps_0_f2h_axi_slave_rvalid),  //                                        .rvalid
		.hps_0_f2h_axi_slave_rready                    (mm_interconnect_1_hps_0_f2h_axi_slave_rready),  //                                        .rready
		.clock_bridge_0_out_clk_clk                    (sys_clk_clk),                                   //                  clock_bridge_0_out_clk.clk
		.mm_bridge_1_reset_reset_bridge_in_reset_reset (sys_rst_reset),                                 // mm_bridge_1_reset_reset_bridge_in_reset.reset
		.mm_bridge_1_m0_address                        (mm_bridge_1_m0_address),                        //                          mm_bridge_1_m0.address
		.mm_bridge_1_m0_waitrequest                    (mm_bridge_1_m0_waitrequest),                    //                                        .waitrequest
		.mm_bridge_1_m0_burstcount                     (mm_bridge_1_m0_burstcount),                     //                                        .burstcount
		.mm_bridge_1_m0_byteenable                     (mm_bridge_1_m0_byteenable),                     //                                        .byteenable
		.mm_bridge_1_m0_read                           (mm_bridge_1_m0_read),                           //                                        .read
		.mm_bridge_1_m0_readdata                       (mm_bridge_1_m0_readdata),                       //                                        .readdata
		.mm_bridge_1_m0_readdatavalid                  (mm_bridge_1_m0_readdatavalid),                  //                                        .readdatavalid
		.mm_bridge_1_m0_write                          (mm_bridge_1_m0_write),                          //                                        .write
		.mm_bridge_1_m0_writedata                      (mm_bridge_1_m0_writedata),                      //                                        .writedata
		.mm_bridge_1_m0_debugaccess                    (mm_bridge_1_m0_debugaccess),                    //                                        .debugaccess
		.mm_bridge_2_m0_address                        (mm_bridge_2_m0_address),                        //                          mm_bridge_2_m0.address
		.mm_bridge_2_m0_waitrequest                    (mm_bridge_2_m0_waitrequest),                    //                                        .waitrequest
		.mm_bridge_2_m0_burstcount                     (mm_bridge_2_m0_burstcount),                     //                                        .burstcount
		.mm_bridge_2_m0_byteenable                     (mm_bridge_2_m0_byteenable),                     //                                        .byteenable
		.mm_bridge_2_m0_read                           (mm_bridge_2_m0_read),                           //                                        .read
		.mm_bridge_2_m0_readdata                       (mm_bridge_2_m0_readdata),                       //                                        .readdata
		.mm_bridge_2_m0_readdatavalid                  (mm_bridge_2_m0_readdatavalid),                  //                                        .readdatavalid
		.mm_bridge_2_m0_write                          (mm_bridge_2_m0_write),                          //                                        .write
		.mm_bridge_2_m0_writedata                      (mm_bridge_2_m0_writedata),                      //                                        .writedata
		.mm_bridge_2_m0_debugaccess                    (mm_bridge_2_m0_debugaccess),                    //                                        .debugaccess
		.mm_bridge_3_m0_address                        (mm_bridge_3_m0_address),                        //                          mm_bridge_3_m0.address
		.mm_bridge_3_m0_waitrequest                    (mm_bridge_3_m0_waitrequest),                    //                                        .waitrequest
		.mm_bridge_3_m0_burstcount                     (mm_bridge_3_m0_burstcount),                     //                                        .burstcount
		.mm_bridge_3_m0_byteenable                     (mm_bridge_3_m0_byteenable),                     //                                        .byteenable
		.mm_bridge_3_m0_read                           (mm_bridge_3_m0_read),                           //                                        .read
		.mm_bridge_3_m0_readdata                       (mm_bridge_3_m0_readdata),                       //                                        .readdata
		.mm_bridge_3_m0_readdatavalid                  (mm_bridge_3_m0_readdatavalid),                  //                                        .readdatavalid
		.mm_bridge_3_m0_write                          (mm_bridge_3_m0_write),                          //                                        .write
		.mm_bridge_3_m0_writedata                      (mm_bridge_3_m0_writedata),                      //                                        .writedata
		.mm_bridge_3_m0_debugaccess                    (mm_bridge_3_m0_debugaccess),                    //                                        .debugaccess
		.mm_bridge_4_m0_address                        (mm_bridge_4_m0_address),                        //                          mm_bridge_4_m0.address
		.mm_bridge_4_m0_waitrequest                    (mm_bridge_4_m0_waitrequest),                    //                                        .waitrequest
		.mm_bridge_4_m0_burstcount                     (mm_bridge_4_m0_burstcount),                     //                                        .burstcount
		.mm_bridge_4_m0_byteenable                     (mm_bridge_4_m0_byteenable),                     //                                        .byteenable
		.mm_bridge_4_m0_read                           (mm_bridge_4_m0_read),                           //                                        .read
		.mm_bridge_4_m0_readdata                       (mm_bridge_4_m0_readdata),                       //                                        .readdata
		.mm_bridge_4_m0_readdatavalid                  (mm_bridge_4_m0_readdatavalid),                  //                                        .readdatavalid
		.mm_bridge_4_m0_write                          (mm_bridge_4_m0_write),                          //                                        .write
		.mm_bridge_4_m0_writedata                      (mm_bridge_4_m0_writedata),                      //                                        .writedata
		.mm_bridge_4_m0_debugaccess                    (mm_bridge_4_m0_debugaccess)                     //                                        .debugaccess
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~hps_0_h2f_reset_reset), // reset_in0.reset
		.clk            (sys_clk_clk),            //       clk.clk
		.reset_out      (sys_rst_reset),          // reset_out.reset
		.reset_req      (),                       // (terminated)
		.reset_req_in0  (1'b0),                   // (terminated)
		.reset_in1      (1'b0),                   // (terminated)
		.reset_req_in1  (1'b0),                   // (terminated)
		.reset_in2      (1'b0),                   // (terminated)
		.reset_req_in2  (1'b0),                   // (terminated)
		.reset_in3      (1'b0),                   // (terminated)
		.reset_req_in3  (1'b0),                   // (terminated)
		.reset_in4      (1'b0),                   // (terminated)
		.reset_req_in4  (1'b0),                   // (terminated)
		.reset_in5      (1'b0),                   // (terminated)
		.reset_req_in5  (1'b0),                   // (terminated)
		.reset_in6      (1'b0),                   // (terminated)
		.reset_req_in6  (1'b0),                   // (terminated)
		.reset_in7      (1'b0),                   // (terminated)
		.reset_req_in7  (1'b0),                   // (terminated)
		.reset_in8      (1'b0),                   // (terminated)
		.reset_req_in8  (1'b0),                   // (terminated)
		.reset_in9      (1'b0),                   // (terminated)
		.reset_req_in9  (1'b0),                   // (terminated)
		.reset_in10     (1'b0),                   // (terminated)
		.reset_req_in10 (1'b0),                   // (terminated)
		.reset_in11     (1'b0),                   // (terminated)
		.reset_req_in11 (1'b0),                   // (terminated)
		.reset_in12     (1'b0),                   // (terminated)
		.reset_req_in12 (1'b0),                   // (terminated)
		.reset_in13     (1'b0),                   // (terminated)
		.reset_req_in13 (1'b0),                   // (terminated)
		.reset_in14     (1'b0),                   // (terminated)
		.reset_req_in14 (1'b0),                   // (terminated)
		.reset_in15     (1'b0),                   // (terminated)
		.reset_req_in15 (1'b0)                    // (terminated)
	);

endmodule
