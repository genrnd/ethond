`define MAX_POS 6 //max word position

`define MAX_POS_L2 4
