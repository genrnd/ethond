`define IP_ETHTYPE         16'h0800 //big endian
`define LOOPBACK_ETHTYPE   16'h9000 //big endian 

`define PTP_ETHTYPE        16'h88F7
`define ARP_ETHTYPE        16'h0806
`define OAM_MAC_ADDRESS    48'h02_00_00_c2_80_01
