`define ICMP_PROTO          8'd1
`define TCP_PROTO           8'd6
`define UDP_PROTO           8'd17

`define SSH_PORT            16'd22  
`define TELNET_PORT         16'd23  
`define ET_DISCOVER_PORT    16'h8018  

`define PTP_EVENT_PORT      16'd319
`define PTP_GENERAL_PORT    16'd320

`define TWAMP_CONTROL_PORT  16'd862


// для DHCP два порта используется
`define DHCP_PORT_A         16'd67
`define DHCP_PORT_B         16'd68

`define DNS_PORT            16'd53

